../chisel/verilog/channel_equalizer.v